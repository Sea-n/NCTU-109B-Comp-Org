`timescale 1ns/1ps

// Author: 0816146 韋詠祥

module ALU(
	src1_i,
	src2_i,
	ctrl_i,
	result_o,
	zero_o
);

// I/O ports
input signed [32-1:0]  src1_i, src2_i;
input [4-1:0] ctrl_i;
output reg [32-1:0] result_o;
output zero_o;

// Parameter

// Main function

endmodule
